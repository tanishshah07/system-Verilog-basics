// driver convert transition lever to pin lever
// monitor coverts opposite
//
//
//steps 
//
//1 -> complete the skeleton first
//2 -> complete and implement the drvier
//3-> completer and implement monitor
//4 -> rest of the fields
//compile it simulate it and make sure that the it will be error free
