`ifndef DEF_SV
`define DEF_SV
parameter SKW_T = 1;
parameter DRAIN_T =20;
typedef enum {IDLE,write,read,simul,res} funct;
`define ADDR_WID 4
`define DEP 16
`define DATA_WID 8 
`endif
