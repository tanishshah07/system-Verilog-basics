
class gen;
int hme;
int x;

endclass

class drv;
gen g1;
task reset();

function new();
 g1=new();
endfunction

endclass

