package pkg;
	
`include "transcation.sv"
`include "generator.sv"
`include "driver.sv"
endpackage
