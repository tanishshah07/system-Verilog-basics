`ifndef INF_SV
`define INF_SV
interface mem_intf(input clk);
logic wr_enb,rd_enb;
//logic [`ADDR_WID-1:0] rd_addr,wr_addr;
//logic [`DATA_WID-1:0] rd_data,wr_data;
logic [3:0] rd_addr,wr_addr;
logic [7:0] rd_data,wr_data;

logic rst=0; //for skeleton zero



//clocking mem_cb@(posedge clk);
  //input 
//endclocking

endinterface
`endif
