`ifndef PKG_SV
`define PKG_SV
//`include "mem_def.sv"
//`include "mem_inter.sv"
package pkg;
event item;
`include "mem_def.sv"
`include "mem_trans.sv"
`include "mem_gen.sv"
`include "mem_driv.sv"
`include "mem_moni.sv"
`include "mem_rfm.sv"
`include "mem_scr.sv"
`include "mem_env.sv"
`include "mem_test.sv"

endpackage
`endif
