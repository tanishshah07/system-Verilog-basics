package pkg;

`include "transcation.sv"
`include "generator.sv"
`include "driver.sv"
`include "and_moni.sv"
`include "ref_mod.sv"
`include "and_scor.sv"
`include "env.sv"
endpackage
