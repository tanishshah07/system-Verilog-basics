////////////////////////////////////////////////
//
//Company_Name : Scaledge
//Author_Name  : TANISH_SHAH
//File_Name    : afifo_driv.sv
//File_Path    : 
//Class_Name   : afifo_driv              
//Project_Name : Asyncronous_FIFO
//Description  :
//
/////////////////////////////////////////////////
`ifndef DRV_SV
`define DRV_SV
class afifo_driv;



endclass
`endif
