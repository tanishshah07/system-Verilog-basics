interface and_intf();
 logic a,b,y;

 modport dut_mp(input a,b,output y);
 
endinterface
