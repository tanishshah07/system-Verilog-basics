class and_transx;
  rand bit a;
  rand bit b;
  bit y;
endclass
