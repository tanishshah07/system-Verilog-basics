`include "intf.sv"
`include "hf.sv"
`include "tb.sv"
module top();
  hf_intf intf();
  hf dut(intf);
  tb test1(intf);
endmodule
