`ifndef DEF_SV
`define DEF_SV

typedef enum {IDLE,write,read} funct;
`define ADDR_WID 4
`define DEP 16
`define DATA_WID 8 

`endif
